interface deserializer_if(input clk);

logic rx_p;
logic rx_n;

endinterface: deserializer_if
