//------------------------------------------------------------
//   Copyright 2010-2018 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//   
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//   
//       http://www.apache.org/licenses/LICENSE-2.0
//   
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------

//
// Class Description:
//
//
class decoder_sequencer extends uvm_sequencer#(decoder_8b10b_trans);

// UVM Factory Registration Macro
//
`uvm_component_utils(decoder_sequencer)

// Standard UVM Methods:
extern function new(string name="decoder_sequencer", 
uvm_component parent = null);

endclass: decoder_sequencer

function decoder_sequencer::new(string name="decoder_sequencer", 
    uvm_component parent = null);
  super.new(name, parent);
endfunction
