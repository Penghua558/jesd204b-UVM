package decoder_8b10b_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
`include "decoder_8b10b_trans.sv"
`include "decoder_8b10b_agent_config.sv"

`include "decoder_8b10b_monitor.sv"
`include "decoder_8b10b_recorder.sv"

`include "decoder_8b10b_agent.sv"
endpackage: decoder_8b10b_agent_pkg
