package apb_agent_dec;
    typedef enum bit {
        WRITE = 1'b1,
        READ = 1'b0
        } op_e;
endpackage: apb_agent_dec
