package enc_bus_dec;
    parameter [7:0] K28_0 = 8'b000_11100;
    parameter [7:0] K28_1 = 8'b001_11100;
    parameter [7:0] K28_2 = 8'b010_11100;
    parameter [7:0] K28_3 = 8'b011_11100;
    parameter [7:0] K28_4 = 8'b100_11100;
    parameter [7:0] K28_5 = 8'b101_11100;
    parameter [7:0] K28_6 = 8'b110_11100;
    parameter [7:0] K28_7 = 8'b111_11100;
    parameter [7:0] K23_7 = 8'b111_10111;
    parameter [7:0] K27_7 = 8'b111_11011;
    parameter [7:0] K29_7 = 8'b111_11101;
    parameter [7:0] K30_7 = 8'b111_11110;
endpackage: enc_bus_dec
