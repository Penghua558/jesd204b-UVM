package deserializer_agent_dec;
    parameter bit[9:0] K_285_MINUS = 10'b001111_1010;
    parameter bit[9:0] K_285_PLUS = 10'b110000_0101;
    bit[9:0] COMMA[2] = {K_285_MINUS, K_285_PLUS};
endpackage: deserializer_agent_dec
