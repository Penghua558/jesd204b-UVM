//------------------------------------------------------------
//   Copyright 2010-2018 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------
package enc_bus_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
`include "enc_bus_trans.sv"
`include "enc_bus_agent_config.sv"

`include "enc_bus_monitor.sv"
`include "enc_bus_driver.sv"
`include "enc_bus_sequencer.sv"
`include "enc_bus_recorder.sv"

`include "enc_bus_agent.sv"

`include "enc_bus_sequences/enc_bus_rand_legal_sequence.sv"
`include "enc_bus_sequences/enc_bus_valid_legal_sequence.sv"
`include "enc_bus_sequences/enc_bus_rand_illegal_sequence.sv"
`include "enc_bus_sequences/enc_bus_valid_illegal_sequence.sv"
endpackage: enc_bus_agent_pkg
