package decoder_8b10b_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
`include "decoder_8b10b_trans.sv"
`include "decoder_8b10b_agent_config.sv"

`include "apb_monitor.sv"
`include "apb_sequencer.sv"
`include "apb_recorder.sv"

`include "apb_agent.sv"

`include "apb_sequences/apb_rand_read_sequence.sv"
`include "apb_sequences/apb_rand_sequence.sv"
endpackage: decoder_8b10b_agent_pkg
