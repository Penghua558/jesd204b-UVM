package cgs2erb_monitor_dec;

typedef bit[7:0] frame_data[];

parameter bit[7:0] R = 8'h1c;

`include "./circular_buffer.svh"

endpackage: cgs2erb_monitor_dec
