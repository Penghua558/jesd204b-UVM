package deserializer_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
`include "deserializer_trans.sv"
`include "decoder_8b10b_agent_config.sv"

`include "decoder_8b10b_monitor.sv"
`include "decoder_8b10b_recorder.sv"

`include "deserializer_agent.sv"
endpackage: deserializer_agent_pkg
