interface decoder_8b10b_if(input clk, input rst_n);

logic [9:0] data;
logic k_error;

endinterface: decoder_8b10b_if
