package deserializer_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
`include "deserializer_trans.sv"
`include "deserializer_agent_config.sv"

`include "deserializer_monitor.sv"
`include "deserializer_recorder.sv"
`include "deserializer_driver.sv"
`include "deserializer_sequencer.sv"

`include "deserializer_agent.sv"
endpackage: deserializer_agent_pkg
