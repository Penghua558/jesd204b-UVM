package table_8b10b_pkg;
    // D word array, value is abcdei, index is EDCBA, running disparity is RD-
    bit [9:0] d_8b_minus[256] = '{
        10'h274,
        10'h1d4,
        10'h2d4,
        10'h31b,
        10'h354,
        10'h29b,
        10'h19b,
        10'h38b,
        10'h394,
        10'h25b,
        10'h15b,
        10'h34b,
        10'hdb ,
        10'h2cb,
        10'h1cb,
        10'h174,
        10'h1b4,
        10'h23b,
        10'h13b,
        10'h32b,
        10'hbb ,
        10'h2ab,
        10'h1ab,
        10'h3a4,
        10'h334,
        10'h26b,
        10'h16b,
        10'h364,
        10'heb ,
        10'h2e4,
        10'h1e4,
        10'h2b4,
        10'h279,
        10'h1d9,
        10'h2d9,
        10'h319,
        10'h359,
        10'h299,
        10'h199,
        10'h389,
        10'h399,
        10'h259,
        10'h159,
        10'h349,
        10'hd9 ,
        10'h2c9,
        10'h1c9,
        10'h179,
        10'h1b9,
        10'h239,
        10'h139,
        10'h329,
        10'hb9 ,
        10'h2a9,
        10'h1a9,
        10'h3a9,
        10'h339,
        10'h269,
        10'h169,
        10'h369,
        10'he9 ,
        10'h2e9,
        10'h1e9,
        10'h2b9,
        10'h275,
        10'h1d5,
        10'h2d5,
        10'h315,
        10'h355,
        10'h295,
        10'h195,
        10'h385,
        10'h395,
        10'h255,
        10'h155,
        10'h345,
        10'hd5 ,
        10'h2c5,
        10'h1c5,
        10'h175,
        10'h1b5,
        10'h235,
        10'h135,
        10'h325,
        10'hb5 ,
        10'h2a5,
        10'h1a5,
        10'h3a5,
        10'h335,
        10'h265,
        10'h165,
        10'h365,
        10'he5 ,
        10'h2e5,
        10'h1e5,
        10'h2b5,
        10'h273,
        10'h1d3,
        10'h2d3,
        10'h31c,
        10'h353,
        10'h29c,
        10'h19c,
        10'h38c,
        10'h393,
        10'h25c,
        10'h15c,
        10'h34c,
        10'hdc ,
        10'h2cc,
        10'h1cc,
        10'h173,
        10'h1b3,
        10'h23c,
        10'h13c,
        10'h32c,
        10'hbc ,
        10'h2ac,
        10'h1ac,
        10'h3a3,
        10'h333,
        10'h26c,
        10'h16c,
        10'h363,
        10'hec ,
        10'h2e3,
        10'h1e3,
        10'h2b3,
        10'h272,
        10'h1d2,
        10'h2d2,
        10'h31d,
        10'h352,
        10'h29d,
        10'h19d,
        10'h38d,
        10'h392,
        10'h25d,
        10'h15d,
        10'h34d,
        10'hdd ,
        10'h2cd,
        10'h1cd,
        10'h172,
        10'h1b2,
        10'h23d,
        10'h13d,
        10'h32d,
        10'hbd ,
        10'h2ad,
        10'h1ad,
        10'h3a2,
        10'h332,
        10'h26d,
        10'h16d,
        10'h362,
        10'hed ,
        10'h2e2,
        10'h1e2,
        10'h2b2,
        10'h27a,
        10'h1da,
        10'h2da,
        10'h31a,
        10'h35a,
        10'h29a,
        10'h19a,
        10'h38a,
        10'h39a,
        10'h25a,
        10'h15a,
        10'h34a,
        10'hda ,
        10'h2ca,
        10'h1ca,
        10'h17a,
        10'h1ba,
        10'h23a,
        10'h13a,
        10'h32a,
        10'hba ,
        10'h2aa,
        10'h1aa,
        10'h3aa,
        10'h33a,
        10'h26a,
        10'h16a,
        10'h36a,
        10'hea ,
        10'h2ea,
        10'h1ea,
        10'h2ba,
        10'h276,
        10'h1d6,
        10'h2d6,
        10'h316,
        10'h356,
        10'h296,
        10'h196,
        10'h386,
        10'h396,
        10'h256,
        10'h156,
        10'h346,
        10'hd6 ,
        10'h2c6,
        10'h1c6,
        10'h176,
        10'h1b6,
        10'h236,
        10'h136,
        10'h326,
        10'hb6 ,
        10'h2a6,
        10'h1a6,
        10'h3a6,
        10'h336,
        10'h266,
        10'h166,
        10'h366,
        10'he6 ,
        10'h2e6,
        10'h1e6,
        10'h2b6,
        10'h271,
        10'h1d1,
        10'h2d1,
        10'h31e,
        10'h351,
        10'h29e,
        10'h19e,
        10'h38e,
        10'h391,
        10'h25e,
        10'h15e,
        10'h34e,
        10'hde ,
        10'h2ce,
        10'h1ce,
        10'h171,
        10'h1b1,
        10'h237,
        10'h137,
        10'h32e,
        10'hb7 ,
        10'h2ae,
        10'h1ae,
        10'h3a1,
        10'h331,
        10'h26e,
        10'h16e,
        10'h361,
        10'hee ,
        10'h2e1,
        10'h1e1,
        10'h2b1
    };

    // D word array, value is abcdei, index is EDCBA, running disparity is RD+
    bit [9:0] d_8b_plus[256] = '{
        10'h18b,
        10'h22b,
        10'h12b,
        10'h314,
        10'hab ,
        10'h294,
        10'h194,
        10'h74 ,
        10'h6b ,
        10'h254,
        10'h154,
        10'h344,
        10'hd4 ,
        10'h2c4,
        10'h1c4,
        10'h28b,
        10'h24b,
        10'h234,
        10'h134,
        10'h324,
        10'hb4 ,
        10'h2a4,
        10'h1a4,
        10'h5b ,
        10'hcb ,
        10'h264,
        10'h164,
        10'h9b ,
        10'he4 ,
        10'h11b,
        10'h21b,
        10'h14b,
        10'h189,
        10'h229,
        10'h129,
        10'h319,
        10'ha9 ,
        10'h299,
        10'h199,
        10'h79 ,
        10'h69 ,
        10'h259,
        10'h159,
        10'h349,
        10'hd9 ,
        10'h2c9,
        10'h1c9,
        10'h289,
        10'h249,
        10'h239,
        10'h139,
        10'h329,
        10'hb9 ,
        10'h2a9,
        10'h1a9,
        10'h59 ,
        10'hc9 ,
        10'h269,
        10'h169,
        10'h99 ,
        10'he9 ,
        10'h119,
        10'h219,
        10'h149,
        10'h185,
        10'h225,
        10'h125,
        10'h315,
        10'ha5 ,
        10'h295,
        10'h195,
        10'h75 ,
        10'h65 ,
        10'h255,
        10'h155,
        10'h345,
        10'hd5 ,
        10'h2c5,
        10'h1c5,
        10'h285,
        10'h245,
        10'h235,
        10'h135,
        10'h325,
        10'hb5 ,
        10'h2a5,
        10'h1a5,
        10'h55 ,
        10'hc5 ,
        10'h265,
        10'h165,
        10'h95 ,
        10'he5 ,
        10'h115,
        10'h215,
        10'h145,
        10'h18c,
        10'h22c,
        10'h12c,
        10'h313,
        10'hac ,
        10'h293,
        10'h193,
        10'h73 ,
        10'h6c ,
        10'h253,
        10'h153,
        10'h343,
        10'hd3 ,
        10'h2c3,
        10'h1c3,
        10'h28c,
        10'h24c,
        10'h233,
        10'h133,
        10'h323,
        10'hb3 ,
        10'h2a3,
        10'h1a3,
        10'h5c ,
        10'hcc ,
        10'h263,
        10'h163,
        10'h9c ,
        10'he3 ,
        10'h11c,
        10'h21c,
        10'h14c,
        10'h18d,
        10'h22d,
        10'h12d,
        10'h312,
        10'had ,
        10'h292,
        10'h192,
        10'h72 ,
        10'h6d ,
        10'h252,
        10'h152,
        10'h342,
        10'hd2 ,
        10'h2c2,
        10'h1c2,
        10'h28d,
        10'h24d,
        10'h232,
        10'h132,
        10'h322,
        10'hb2 ,
        10'h2a2,
        10'h1a2,
        10'h5d ,
        10'hcd ,
        10'h262,
        10'h162,
        10'h9d ,
        10'he2 ,
        10'h11d,
        10'h21d,
        10'h14d,
        10'h18a,
        10'h22a,
        10'h12a,
        10'h31a,
        10'haa ,
        10'h29a,
        10'h19a,
        10'h7a ,
        10'h6a ,
        10'h25a,
        10'h15a,
        10'h34a,
        10'hda ,
        10'h2ca,
        10'h1ca,
        10'h28a,
        10'h24a,
        10'h23a,
        10'h13a,
        10'h32a,
        10'hba ,
        10'h2aa,
        10'h1aa,
        10'h5a ,
        10'hca ,
        10'h26a,
        10'h16a,
        10'h9a ,
        10'hea ,
        10'h11a,
        10'h21a,
        10'h14a,
        10'h186,
        10'h226,
        10'h126,
        10'h316,
        10'ha6 ,
        10'h296,
        10'h196,
        10'h76 ,
        10'h66 ,
        10'h256,
        10'h156,
        10'h346,
        10'hd6 ,
        10'h2c6,
        10'h1c6,
        10'h286,
        10'h246,
        10'h236,
        10'h136,
        10'h326,
        10'hb6 ,
        10'h2a6,
        10'h1a6,
        10'h56 ,
        10'hc6 ,
        10'h266,
        10'h166,
        10'h96 ,
        10'he6 ,
        10'h116,
        10'h216,
        10'h146,
        10'h18e,
        10'h22e,
        10'h12e,
        10'h311,
        10'hae ,
        10'h291,
        10'h191,
        10'h71 ,
        10'h6e ,
        10'h251,
        10'h151,
        10'h348,
        10'hd1 ,
        10'h2c8,
        10'h1c8,
        10'h28e,
        10'h24e,
        10'h231,
        10'h131,
        10'h321,
        10'hb1 ,
        10'h2a1,
        10'h1a1,
        10'h5e ,
        10'hce ,
        10'h261,
        10'h161,
        10'h9e ,
        10'he1 ,
        10'h11e,
        10'h21e,
        10'h14e
        };


    // K word array, value is abcdeifghj, index is HGFEDCBA, running disparity
    // is RD-
    bit [9:0] k_8b_minus[byte] = '{
        8'b000_11100:10'b001111_0100,
        8'b001_11100:10'b001111_1001,
        8'b010_11100:10'b001111_0101,
        8'b011_11100:10'b001111_0011,
        8'b100_11100:10'b001111_0010,
        8'b101_11100:10'b001111_1010,
        8'b110_11100:10'b001111_0110,
        8'b111_11100:10'b001111_1000,
        8'b111_10111:10'b111010_1000,
        8'b111_11011:10'b110110_1000,
        8'b111_11101:10'b101110_1000,
        8'b111_11110:10'b011110_1000
    };

    // K word array, value is abcdeifghj, index is HGFEDCBA, running disparity
    // is RD+
    bit [9:0] k_8b_plus[byte] = '{
        8'b000_11100:10'b110000_1011,
        8'b001_11100:10'b110000_0110,
        8'b010_11100:10'b110000_1010,
        8'b011_11100:10'b110000_1100,
        8'b100_11100:10'b110000_1101,
        8'b101_11100:10'b110000_0101,
        8'b110_11100:10'b110000_1001,
        8'b111_11100:10'b110000_0111,
        8'b111_10111:10'b000101_0111,
        8'b111_11011:10'b001001_0111,
        8'b111_11101:10'b010001_0111,
        8'b111_11110:10'b100001_0111
    };
endpackage: table_8b10b_pkg
