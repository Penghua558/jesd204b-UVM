interface deserializer_if(input bitclk, input device_clk, input rst_n);
logic rx_p;
logic rx_n;
logic sync_n;

endinterface: deserializer_if
