interface enc_bus_if(input clk, input rst_n);

// HGFEDCBA
logic [7:0] data;
logic valid;
logic k;

endinterface: enc_bus_if
